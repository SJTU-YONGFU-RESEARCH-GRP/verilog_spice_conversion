* Standard Cell Library SPICE Models
* Generic technology library for ngspice
* Uses generic MOSFET models - replace with technology-specific models as needed
*
* Note: This library requires MOSFET model definitions. Include the technology
* model file in your main SPICE netlist:

* ============================================================================
* Generic 0.18um CMOS Technology Models
* ============================================================================

* NMOS Transistor Model
* Level 1 (Shichman-Hodges) model with generic 0.18um CMOS parameters
.model NMOS NMOS (LEVEL=1 VTO=0.7 KP=200u GAMMA=0.5 PHI=0.7 LAMBDA=0.05 TOX=4.1n NSUB=1e17 LD=0.08u WD=0.08u UO=350 CJ=0.0004 CJSW=5e-10 PB=0.9 MJ=0.5 MJSW=0.3 RD=0 RS=0 RSH=0 IS=1e-15 JS=0 N=1 TPG=1 XJ=0 CGSO=0 CGDO=0 CGBO=0)

* PMOS Transistor Model
* Level 1 (Shichman-Hodges) model with generic 0.18um CMOS parameters
.model PMOS PMOS (LEVEL=1 VTO=-0.7 KP=100u GAMMA=0.5 PHI=0.7 LAMBDA=0.05 TOX=4.1n NSUB=1e17 LD=0.08u WD=0.08u UO=100 CJ=0.0004 CJSW=5e-10 PB=0.9 MJ=0.5 MJSW=0.3 RD=0 RS=0 RSH=0 IS=1e-15 JS=0 N=1 TPG=1 XJ=0 CGSO=0 CGDO=0 CGBO=0)

* ============================================================================
* Basic Gates
* ============================================================================

* Inverter
* CMOS inverter: PMOS pull-up, NMOS pull-down
.SUBCKT INV A Y
* PMOS: source=VDD, drain=Y, gate=A, bulk=VDD
M1 Y A VDD VDD PMOS W=2u L=0.18u
* NMOS: source=VSS, drain=Y, gate=A, bulk=VSS
M2 Y A VSS VSS NMOS W=1u L=0.18u
.ENDS INV

* Buffer
* Two inverters in series for signal buffering
.SUBCKT BUF A Y
X1 A Y_int INV
X2 Y_int Y INV
.ENDS BUF

* ============================================================================
* 2-Input Gates
* ============================================================================

* 2-input NAND
* CMOS NAND: parallel PMOS pull-up, series NMOS pull-down
.SUBCKT NAND2 A B Y
* PMOS pull-up network (parallel)
M1 Y A VDD VDD PMOS W=2u L=0.18u
M2 Y B VDD VDD PMOS W=2u L=0.18u
* NMOS pull-down network (series)
M3 Y A net1 VSS NMOS W=1u L=0.18u
M4 net1 B VSS VSS NMOS W=1u L=0.18u
.ENDS NAND2

* 2-input NOR
* CMOS NOR: series PMOS pull-up, parallel NMOS pull-down
.SUBCKT NOR2 A B Y
* PMOS pull-up network (series)
M1 Y A net1 VDD PMOS W=2u L=0.18u
M2 net1 B VDD VDD PMOS W=2u L=0.18u
* NMOS pull-down network (parallel)
M3 Y A VSS VSS NMOS W=1u L=0.18u
M4 Y B VSS VSS NMOS W=1u L=0.18u
.ENDS NOR2

* 2-input AND
* AND = NAND + INV
.SUBCKT AND2 A B Y
X1 A B Y_int NAND2
X2 Y_int Y INV
.ENDS AND2

* 2-input OR
* OR = NOR + INV
.SUBCKT OR2 A B Y
X1 A B Y_int NOR2
X2 Y_int Y INV
.ENDS OR2

* 2-input XOR
* CMOS XOR implementation using standard logic gates
* XOR = (A & !B) | (!A & B) = (A | B) & (!A | !B)
.SUBCKT XOR2 A B Y
* Generate complements
X1 A A_bar INV
X2 B B_bar INV
* Intermediate signals: (A & B_bar) and (A_bar & B)
X3 A B_bar n1 AND2
X4 A_bar B n2 AND2
* OR the intermediate signals
X5 n1 n2 Y OR2
.ENDS XOR2

* 2-input XNOR
* XNOR = XOR + INV
.SUBCKT XNOR2 A B Y
X1 A B Y_int XOR2
X2 Y_int Y INV
.ENDS XNOR2

* ============================================================================
* 3-Input Gates
* ============================================================================

* 3-input NAND
* CMOS NAND: parallel PMOS pull-up, series NMOS pull-down
.SUBCKT NAND3 A B C Y
* PMOS pull-up network (parallel)
M1 Y A VDD VDD PMOS W=2u L=0.18u
M2 Y B VDD VDD PMOS W=2u L=0.18u
M3 Y C VDD VDD PMOS W=2u L=0.18u
* NMOS pull-down network (series)
M4 Y A net1 VSS NMOS W=1u L=0.18u
M5 net1 B net2 VSS NMOS W=1u L=0.18u
M6 net2 C VSS VSS NMOS W=1u L=0.18u
.ENDS NAND3

* 3-input NOR
* CMOS NOR: series PMOS pull-up, parallel NMOS pull-down
.SUBCKT NOR3 A B C Y
* PMOS pull-up network (series)
M1 Y A net1 VDD PMOS W=2u L=0.18u
M2 net1 B net2 VDD PMOS W=2u L=0.18u
M3 net2 C VDD VDD PMOS W=2u L=0.18u
* NMOS pull-down network (parallel)
M4 Y A VSS VSS NMOS W=1u L=0.18u
M5 Y B VSS VSS NMOS W=1u L=0.18u
M6 Y C VSS VSS NMOS W=1u L=0.18u
.ENDS NOR3

* ============================================================================
* Sequential Elements
* ============================================================================

* D Flip-Flop (Master-Slave)
* Master-slave D flip-flop using transmission gates
.SUBCKT DFF D CLK Q QN
* Generate clock and clock bar
X1 CLK CLK_bar INV
* Master latch (transparent when CLK=0)
X2 D CLK CLK_bar master_out TGATE
X3 master_out master_q INV
X4 master_q master_out INV
* Slave latch (transparent when CLK=1)
X5 master_q CLK_bar CLK slave_out TGATE
X6 slave_out QN INV
X7 QN Q INV
.ENDS DFF

* D Flip-Flop with Reset
* Master-slave D flip-flop with asynchronous reset
.SUBCKT DFFR D CLK RST Q QN
* Generate clock and clock bar
X1 CLK CLK_bar INV
* Reset logic: when RST=1, force Q=0
X2 RST D net1 NOR2
X3 net1 CLK CLK_bar master_out TGATE
X4 master_out master_q INV
X5 master_q master_out INV
* Slave latch with reset
X6 master_q CLK_bar CLK slave_out TGATE
X7 RST slave_out QN NOR2
X8 QN Q INV
.ENDS DFFR

* ============================================================================
* Helper Subcircuits
* ============================================================================

* Transmission Gate (for use in sequential elements)
* Complementary pass gate: passes signal when EN=1, EN_bar=0
.SUBCKT TGATE IN OUT EN EN_bar
* PMOS pass transistor (active when EN_bar=0, i.e., EN=1)
M1 OUT EN_bar IN VDD PMOS W=2u L=0.18u
* NMOS pass transistor (active when EN=1)
M2 OUT EN IN VSS NMOS W=1u L=0.18u
.ENDS TGATE
